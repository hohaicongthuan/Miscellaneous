module featuremap4(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.053731956),
	.w1(0.10092049),
	.w2(-0.09923359),
	.w3(0.0058972454),
	.w4(-0.014974821),
	.w5(0.08036631),
	.w6(-0.08273384),
	.w7(-0.0425488),
	.w8(-0.055765543),
	.w9(0.065507315),
	.w10(0.04099769),
	.w11(0.015825808),
	.w12(-0.08832933),
	.w13(-0.012153113),
	.w14(-0.10947188),
	.w15(-0.09480668),
	.w16(0.08207682),
	.w17(-0.05715896),
	.w18(0.07945019),
	.w19(-0.06776747),
	.w20(0.06566027),
	.w21(-0.081792995),
	.w22(0.08097058),
	.w23(-0.009838002),
	.w24(0.0433402),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.07032161),
	.w1(-0.09053616),
	.w2(0.045173693),
	.w3(0.067935474),
	.w4(-0.073682405),
	.w5(0.060056332),
	.w6(-0.07589911),
	.w7(0.106547676),
	.w8(0.0022574768),
	.w9(-0.0816233),
	.w10(-0.02951384),
	.w11(-0.08103216),
	.w12(0.032579437),
	.w13(-0.041619767),
	.w14(-0.06459623),
	.w15(-0.09769),
	.w16(0.037186313),
	.w17(-0.028580483),
	.w18(0.057503924),
	.w19(-0.044959716),
	.w20(-0.017739804),
	.w21(-0.048362505),
	.w22(-0.011113269),
	.w23(-0.033565227),
	.w24(0.09422937),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.10517619),
	.w1(-0.06281464),
	.w2(-0.104100436),
	.w3(0.0015249532),
	.w4(-0.08494289),
	.w5(-0.08417986),
	.w6(0.1029205),
	.w7(0.09960193),
	.w8(-0.10759574),
	.w9(-0.034404345),
	.w10(-0.10309433),
	.w11(-0.1127541),
	.w12(-0.11468618),
	.w13(-0.073209986),
	.w14(0.020000048),
	.w15(-0.11433289),
	.w16(-0.07476218),
	.w17(0.025880555),
	.w18(0.041168228),
	.w19(-0.032675326),
	.w20(0.09212787),
	.w21(-0.063891746),
	.w22(-0.1058366),
	.w23(0.06992726),
	.w24(0.094000675),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule