Ring Oscillator
.include 45nm_LP.lib SS
.option TEMP = -40C

// Capacitance value for Ring Oscillator
.param cap_val = 1p
// Resistance value for Ring Oscillator
.param res_val = 1k

    * Syntax for MOSFET
    * MXXXXXXX nd ng ns nb mname <m = val > <l = val> <w = val>

    // Pull-down network
    M1 gate_1_out RgOsc_Out 0 0 NMOS
    M2 gate_2_out res_1_out 0 0 NMOS
    M3 gate_3_out res_2_out 0 0 NMOS

    // Pull-up network
    M4 gate_1_out RgOsc_Out vdd vdd PMOS
    M5 gate_2_out res_1_out vdd vdd PMOS
    M6 gate_3_out res_2_out vdd vdd PMOS

    // Resistors
    R1 gate_1_out res_1_out res_val
    R2 gate_2_out res_2_out res_val
    R3 gate_3_out RgOsc_Out res_val

    // Capacitors
    C1 res_1_out 0 cap_val
    C2 res_2_out 0 cap_val
    C3 RgOsc_Out 0 cap_val

    // Power
    V1 vdd 0 dc 0.9V

.control
    * General form: .tran tstep tstop <tstart<tmax>> <uic>
    tran 1ns 5us
    plot RgOsc_Out
.endc

.end