module featuremap12(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.047969095),
	.w1(0.032378945),
	.w2(-0.030710788),
	.w3(-0.078425445),
	.w4(-0.011341424),
	.w5(0.060580853),
	.w6(-0.08134082),
	.w7(-0.06265078),
	.w8(0.011671211),
	.w9(0.045993235),
	.w10(0.07268335),
	.w11(0.06013741),
	.w12(0.06410545),
	.w13(0.07586355),
	.w14(-0.0736486),
	.w15(-0.0056753983),
	.w16(-0.021568032),
	.w17(-0.08066696),
	.w18(0.029507857),
	.w19(-0.034028728),
	.w20(0.05459459),
	.w21(0.07559184),
	.w22(0.061054666),
	.w23(-0.076866716),
	.w24(0.019986326),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.024601767),
	.w1(-0.065144435),
	.w2(0.007193497),
	.w3(-0.054081768),
	.w4(0.07131391),
	.w5(0.060041614),
	.w6(-0.012358125),
	.w7(0.07198363),
	.w8(0.035235535),
	.w9(-0.03526739),
	.w10(0.05396529),
	.w11(0.06885519),
	.w12(-0.044902276),
	.w13(0.00016314149),
	.w14(-0.06755858),
	.w15(-0.02742384),
	.w16(0.04014766),
	.w17(-0.0732805),
	.w18(0.06983314),
	.w19(0.050552662),
	.w20(-0.072142065),
	.w21(0.016759666),
	.w22(0.012828395),
	.w23(0.06787535),
	.w24(0.009292864),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.025029764),
	.w1(0.055211853),
	.w2(-0.061844707),
	.w3(0.015639167),
	.w4(-0.07641208),
	.w5(0.0655352),
	.w6(-0.024773786),
	.w7(0.07238955),
	.w8(-0.06723982),
	.w9(0.06967114),
	.w10(-0.073524475),
	.w11(-0.0697196),
	.w12(0.014829932),
	.w13(0.0031695643),
	.w14(-0.011412634),
	.w15(-0.06653436),
	.w16(-0.0155703705),
	.w17(-0.023305064),
	.w18(0.024162956),
	.w19(0.024803258),
	.w20(0.004762873),
	.w21(0.07774216),
	.w22(-0.009455695),
	.w23(-0.02698607),
	.w24(0.022266345),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.077563725),
	.w1(-0.02029397),
	.w2(-0.0437259),
	.w3(0.009887468),
	.w4(-0.06975821),
	.w5(0.057082914),
	.w6(0.07493016),
	.w7(0.043465316),
	.w8(0.0528926),
	.w9(0.05021944),
	.w10(0.045034584),
	.w11(-0.0695652),
	.w12(-0.04106879),
	.w13(0.075607635),
	.w14(0.050028693),
	.w15(0.043868337),
	.w16(-0.037978873),
	.w17(0.037530564),
	.w18(0.0684016),
	.w19(-0.071496),
	.w20(-0.008254097),
	.w21(-0.061833855),
	.w22(-0.027162867),
	.w23(0.021607257),
	.w24(-0.07630138),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.025554841),
	.w1(-0.037857495),
	.w2(-0.02679258),
	.w3(0.0250949),
	.w4(-0.067611754),
	.w5(-0.040479157),
	.w6(0.021644974),
	.w7(-0.004700307),
	.w8(0.07117165),
	.w9(0.023271007),
	.w10(-0.05494548),
	.w11(0.060320836),
	.w12(0.021241087),
	.w13(-0.030658811),
	.w14(-0.042580783),
	.w15(-0.06711792),
	.w16(-0.01767439),
	.w17(0.028664205),
	.w18(0.03383597),
	.w19(-0.010121118),
	.w20(-0.06401369),
	.w21(-0.04409056),
	.w22(0.045740392),
	.w23(0.051946223),
	.w24(-0.026693514),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.0011130627),
	.w1(0.046686135),
	.w2(0.074049324),
	.w3(-0.020362921),
	.w4(-0.012623156),
	.w5(-0.014877567),
	.w6(0.037026208),
	.w7(0.018364606),
	.w8(0.060956925),
	.w9(-0.046597153),
	.w10(0.016872777),
	.w11(-0.040854305),
	.w12(0.03518262),
	.w13(0.042681076),
	.w14(-0.036554974),
	.w15(-0.074818924),
	.w16(-0.013042277),
	.w17(0.0026968715),
	.w18(-0.041752256),
	.w19(0.030116087),
	.w20(-0.040027365),
	.w21(-0.030106734),
	.w22(-0.05924221),
	.w23(-0.04496097),
	.w24(0.03301918),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule