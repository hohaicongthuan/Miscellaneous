module featuremap14(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.048569363),
	.w1(-0.055602904),
	.w2(0.021932354),
	.w3(0.07805265),
	.w4(-0.05487108),
	.w5(-0.029242262),
	.w6(-0.030690495),
	.w7(0.06074675),
	.w8(-0.055720445),
	.w9(0.08142041),
	.w10(0.019076098),
	.w11(0.0690419),
	.w12(-0.06044546),
	.w13(0.064893425),
	.w14(0.022733072),
	.w15(0.010568406),
	.w16(-0.025863197),
	.w17(-0.030991646),
	.w18(0.035909183),
	.w19(0.039055962),
	.w20(-0.021843692),
	.w21(-0.046563186),
	.w22(-0.047251042),
	.w23(0.048582204),
	.w24(0.025325757),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.045152728),
	.w1(0.050620776),
	.w2(0.078305244),
	.w3(0.063854925),
	.w4(0.037190028),
	.w5(0.044129953),
	.w6(0.011970377),
	.w7(0.003521884),
	.w8(0.027989272),
	.w9(0.059175253),
	.w10(0.04547186),
	.w11(0.011461349),
	.w12(-0.068958946),
	.w13(-0.070861876),
	.w14(-0.0573405),
	.w15(0.04594458),
	.w16(-0.047596455),
	.w17(0.027119145),
	.w18(-0.053870942),
	.w19(-0.023766048),
	.w20(-0.03923816),
	.w21(-0.02128883),
	.w22(-0.05350155),
	.w23(-0.0658499),
	.w24(-0.04831147),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.023072962),
	.w1(0.023432104),
	.w2(0.06306894),
	.w3(0.047719095),
	.w4(0.06071501),
	.w5(0.057582345),
	.w6(-0.03617429),
	.w7(0.07883309),
	.w8(-0.06786697),
	.w9(0.072177514),
	.w10(0.022713196),
	.w11(-0.06416801),
	.w12(-0.027329192),
	.w13(-0.004996951),
	.w14(-0.04438495),
	.w15(-0.024607413),
	.w16(0.023619132),
	.w17(-0.029082986),
	.w18(0.033643607),
	.w19(-0.048601836),
	.w20(-0.028792433),
	.w21(-0.06709368),
	.w22(0.042630434),
	.w23(0.028666444),
	.w24(0.025979111),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.062948614),
	.w1(0.020439932),
	.w2(-0.06960113),
	.w3(0.075500354),
	.w4(0.024018776),
	.w5(-0.061415464),
	.w6(0.010021341),
	.w7(-0.048368312),
	.w8(-0.038776904),
	.w9(0.07597877),
	.w10(0.07586495),
	.w11(-0.008967136),
	.w12(0.060843218),
	.w13(-0.058437124),
	.w14(-0.06549418),
	.w15(0.0009963983),
	.w16(-0.04045256),
	.w17(0.080736026),
	.w18(-0.0629337),
	.w19(0.06714359),
	.w20(-0.019849844),
	.w21(0.033223078),
	.w22(-0.052087706),
	.w23(0.038313836),
	.w24(0.08155424),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.050758727),
	.w1(-0.06109656),
	.w2(0.064647585),
	.w3(0.033457097),
	.w4(0.012055232),
	.w5(-0.075036675),
	.w6(-0.055352286),
	.w7(0.0116621),
	.w8(0.013595931),
	.w9(0.036040116),
	.w10(-0.04085882),
	.w11(0.010664359),
	.w12(-0.03413021),
	.w13(0.06357397),
	.w14(0.023849268),
	.w15(0.04949363),
	.w16(0.07143774),
	.w17(-0.0659436),
	.w18(-0.07630439),
	.w19(-0.011498832),
	.w20(0.0119317835),
	.w21(0.071251966),
	.w22(-0.00286524),
	.w23(0.027346129),
	.w24(-0.03881536),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.068387195),
	.w1(-0.07152066),
	.w2(-0.049409524),
	.w3(-0.042023215),
	.w4(0.037305936),
	.w5(-0.028131165),
	.w6(0.06603735),
	.w7(0.014955862),
	.w8(0.03215941),
	.w9(-0.034549583),
	.w10(0.07119342),
	.w11(-0.03625615),
	.w12(0.07097673),
	.w13(-0.0692129),
	.w14(-0.049184214),
	.w15(0.029040566),
	.w16(-0.07839479),
	.w17(-0.03164348),
	.w18(-0.03927546),
	.w19(0.017905433),
	.w20(-0.041415833),
	.w21(0.022773825),
	.w22(0.03236646),
	.w23(-0.08109808),
	.w24(0.0065435786),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule