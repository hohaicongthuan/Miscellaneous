module featuremap2(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.030423341),
	.w1(-0.056152344),
	.w2(-0.06998253),
	.w3(-0.010521508),
	.w4(-0.010235056),
	.w5(0.0074314624),
	.w6(-0.059371848),
	.w7(0.053534314),
	.w8(0.0063912887),
	.w9(-0.024525793),
	.w10(0.074516974),
	.w11(-0.013883593),
	.w12(-0.020458963),
	.w13(0.033723608),
	.w14(0.038230468),
	.w15(-0.015556232),
	.w16(-0.04266057),
	.w17(-0.007147764),
	.w18(-0.08296057),
	.w19(-0.08161277),
	.w20(-0.028225081),
	.w21(0.104730904),
	.w22(0.034109417),
	.w23(-0.058339424),
	.w24(-0.014371923),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.020120464),
	.w1(-0.053495966),
	.w2(0.00075801666),
	.w3(-0.063529655),
	.w4(-0.10728907),
	.w5(0.07800893),
	.w6(0.070428364),
	.w7(0.08460615),
	.w8(0.015466731),
	.w9(-0.0030689985),
	.w10(-0.026199395),
	.w11(-0.041891117),
	.w12(-0.038862094),
	.w13(-0.042934965),
	.w14(-0.048882827),
	.w15(0.0055697183),
	.w16(-0.05071229),
	.w17(0.0038303325),
	.w18(0.03102156),
	.w19(-0.093849786),
	.w20(-0.08581161),
	.w21(-0.024129083),
	.w22(0.014517187),
	.w23(0.06441791),
	.w24(-0.11281344),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07076335),
	.w1(-0.11308664),
	.w2(0.06587821),
	.w3(0.073534004),
	.w4(0.11332264),
	.w5(0.090997815),
	.w6(-0.08115148),
	.w7(0.048805658),
	.w8(0.047300376),
	.w9(-0.10739313),
	.w10(0.030421373),
	.w11(-0.022809932),
	.w12(0.023424461),
	.w13(-0.05407454),
	.w14(-0.10518278),
	.w15(-0.11202605),
	.w16(-0.051768214),
	.w17(0.07515378),
	.w18(-0.0013588358),
	.w19(0.020855052),
	.w20(-0.075723045),
	.w21(-0.0582456),
	.w22(0.10747288),
	.w23(0.09061136),
	.w24(-0.022027208),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule