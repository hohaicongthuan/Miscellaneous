module featuremap3(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.049541157),
	.w1(-0.036977723),
	.w2(-0.039385602),
	.w3(0.047036443),
	.w4(0.04333655),
	.w5(0.04525786),
	.w6(-0.013537045),
	.w7(0.05034963),
	.w8(-0.028000437),
	.w9(0.048418477),
	.w10(0.07211699),
	.w11(-0.067041844),
	.w12(0.032285955),
	.w13(-0.015241966),
	.w14(0.03260673),
	.w15(0.00848289),
	.w16(-0.014118469),
	.w17(-0.008890087),
	.w18(-0.06648441),
	.w19(0.07969507),
	.w20(-0.050741225),
	.w21(0.04908321),
	.w22(-0.061721347),
	.w23(0.05866457),
	.w24(0.004245017),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07884243),
	.w1(0.054829564),
	.w2(-0.037117302),
	.w3(0.055733144),
	.w4(0.01027402),
	.w5(0.040466115),
	.w6(0.04292336),
	.w7(0.007801591),
	.w8(0.040651936),
	.w9(0.054280475),
	.w10(0.0036152273),
	.w11(0.05345053),
	.w12(-0.01049236),
	.w13(2.3360155e-07),
	.w14(0.015805997),
	.w15(0.039522793),
	.w16(0.056724444),
	.w17(0.027126465),
	.w18(0.045827992),
	.w19(0.04841101),
	.w20(-0.026320277),
	.w21(-0.051111475),
	.w22(0.08068999),
	.w23(-0.021355368),
	.w24(-0.05070907),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.04498183),
	.w1(0.052545067),
	.w2(-0.004693386),
	.w3(0.015602326),
	.w4(-0.014585604),
	.w5(-0.0041847187),
	.w6(0.016754605),
	.w7(-0.049548086),
	.w8(-0.057535905),
	.w9(-0.065861925),
	.w10(0.030443188),
	.w11(0.031122403),
	.w12(-0.02970714),
	.w13(0.07989688),
	.w14(-0.017415024),
	.w15(-0.026667817),
	.w16(0.0784851),
	.w17(-0.07465886),
	.w18(0.010085698),
	.w19(0.004321736),
	.w20(0.07528085),
	.w21(-0.029840827),
	.w22(-0.025038242),
	.w23(-0.05420619),
	.w24(0.036789693),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.05757409),
	.w1(-0.052286968),
	.w2(0.07083103),
	.w3(0.033827323),
	.w4(0.0016376929),
	.w5(0.053794242),
	.w6(0.01515568),
	.w7(0.07414045),
	.w8(-0.008679397),
	.w9(-0.05875633),
	.w10(-0.06964188),
	.w11(-0.010421481),
	.w12(0.012448967),
	.w13(0.0659304),
	.w14(0.0020538736),
	.w15(-0.068027146),
	.w16(0.07493238),
	.w17(-0.028651794),
	.w18(-0.014126635),
	.w19(0.043376304),
	.w20(0.0450161),
	.w21(-0.0644084),
	.w22(0.034790356),
	.w23(-0.024261585),
	.w24(0.029639238),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.06143745),
	.w1(-0.06598046),
	.w2(0.03973323),
	.w3(0.009966503),
	.w4(0.069966525),
	.w5(-0.07183635),
	.w6(0.04308797),
	.w7(-0.07612876),
	.w8(0.069509424),
	.w9(-0.036853917),
	.w10(0.032642625),
	.w11(-0.076561354),
	.w12(-0.05687969),
	.w13(0.03539673),
	.w14(0.0487948),
	.w15(-0.06512963),
	.w16(0.0701495),
	.w17(0.0112812035),
	.w18(-0.01718011),
	.w19(0.01978576),
	.w20(-0.03520288),
	.w21(-0.023493892),
	.w22(-0.007637077),
	.w23(-0.006292087),
	.w24(0.034936532),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.0069389394),
	.w1(0.06596355),
	.w2(-0.03112478),
	.w3(0.022277616),
	.w4(-0.063071094),
	.w5(0.07667785),
	.w6(0.07544057),
	.w7(-0.028869813),
	.w8(0.08161618),
	.w9(0.013638019),
	.w10(-0.06319652),
	.w11(0.005963984),
	.w12(-0.02310919),
	.w13(-0.052282423),
	.w14(0.05685528),
	.w15(-0.035416145),
	.w16(0.022647291),
	.w17(0.037967786),
	.w18(-0.026850007),
	.w19(0.0780895),
	.w20(0.020250052),
	.w21(0.06151888),
	.w22(-0.0775723),
	.w23(-0.032157347),
	.w24(-0.07791771),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule