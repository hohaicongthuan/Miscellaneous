module featuremap15(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.009665956),
	.w1(-0.039327357),
	.w2(0.06688603),
	.w3(-0.0431305),
	.w4(-0.043725003),
	.w5(-0.069012),
	.w6(0.00079464435),
	.w7(0.06575749),
	.w8(0.0436148),
	.w9(-0.055099502),
	.w10(-0.007815763),
	.w11(-0.03260188),
	.w12(0.0106954565),
	.w13(-0.032576058),
	.w14(0.07542021),
	.w15(-0.013485681),
	.w16(0.0140547445),
	.w17(-0.07190136),
	.w18(-0.0135741),
	.w19(0.070923105),
	.w20(-0.034659542),
	.w21(0.0520814),
	.w22(-0.052374434),
	.w23(0.035859436),
	.w24(-0.01693366),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.046551485),
	.w1(0.034470517),
	.w2(-0.07904915),
	.w3(0.009045227),
	.w4(0.05307328),
	.w5(-0.054638118),
	.w6(0.019321933),
	.w7(-0.016877342),
	.w8(-0.0612412),
	.w9(-0.067305855),
	.w10(-0.010246261),
	.w11(0.0034575074),
	.w12(-0.06806911),
	.w13(-0.054544903),
	.w14(-0.048440963),
	.w15(-0.035168197),
	.w16(-0.035695195),
	.w17(0.013377972),
	.w18(-0.05957553),
	.w19(-0.04715815),
	.w20(-0.07437061),
	.w21(0.012847151),
	.w22(-0.046133745),
	.w23(-0.02318765),
	.w24(-0.024006726),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.051763758),
	.w1(0.08046655),
	.w2(-0.058650896),
	.w3(0.065408826),
	.w4(-0.032456756),
	.w5(0.015235552),
	.w6(-0.015102905),
	.w7(0.07655514),
	.w8(0.041911777),
	.w9(-0.009496565),
	.w10(0.06649287),
	.w11(0.018750798),
	.w12(0.022921432),
	.w13(0.07354074),
	.w14(-0.044896066),
	.w15(0.012944378),
	.w16(0.0130197145),
	.w17(0.07747907),
	.w18(-0.025418332),
	.w19(-0.0019144036),
	.w20(-0.050064366),
	.w21(-0.0280164),
	.w22(-0.008943163),
	.w23(0.04849729),
	.w24(0.039165724),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.024149494),
	.w1(-0.009486452),
	.w2(-0.02670788),
	.w3(-0.06553024),
	.w4(-0.07140924),
	.w5(-0.022103779),
	.w6(0.0027072474),
	.w7(-0.042716283),
	.w8(-0.017579937),
	.w9(-0.01665798),
	.w10(-0.08162123),
	.w11(-0.01032951),
	.w12(0.0074460786),
	.w13(0.04591381),
	.w14(-0.040205114),
	.w15(-0.05385673),
	.w16(0.0038555644),
	.w17(-0.010814029),
	.w18(0.04420156),
	.w19(-0.052601445),
	.w20(-0.0435204),
	.w21(0.019889878),
	.w22(-0.024490582),
	.w23(-0.0064130244),
	.w24(0.011068704),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.032775067),
	.w1(0.049033046),
	.w2(-0.05460663),
	.w3(0.028892638),
	.w4(-0.02638992),
	.w5(-0.002921197),
	.w6(0.043691892),
	.w7(0.017364314),
	.w8(0.01932314),
	.w9(-0.017123578),
	.w10(0.034007635),
	.w11(0.07084853),
	.w12(-0.08071704),
	.w13(0.07433321),
	.w14(-0.06362025),
	.w15(0.065267965),
	.w16(0.025292352),
	.w17(-0.005525368),
	.w18(-0.055117693),
	.w19(0.0018965721),
	.w20(-0.045194115),
	.w21(-0.004476954),
	.w22(0.0041975863),
	.w23(0.07206266),
	.w24(0.049665414),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.03037486),
	.w1(0.03311778),
	.w2(0.037853293),
	.w3(-0.026783187),
	.w4(-0.03833163),
	.w5(0.041255455),
	.w6(0.016607387),
	.w7(-0.01811649),
	.w8(0.008709843),
	.w9(0.07151776),
	.w10(0.05988805),
	.w11(-0.053598113),
	.w12(0.073628195),
	.w13(0.030062573),
	.w14(-0.018366707),
	.w15(0.024257166),
	.w16(-0.036632236),
	.w17(-0.059739772),
	.w18(0.023942145),
	.w19(0.075425096),
	.w20(-0.053787168),
	.w21(-0.07192028),
	.w22(0.015140135),
	.w23(0.075386606),
	.w24(0.06710169),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule