module featuremap5(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.06940607),
	.w1(0.023634832),
	.w2(0.040496524),
	.w3(0.0070020217),
	.w4(-0.06493699),
	.w5(0.04570214),
	.w6(-0.015007771),
	.w7(-0.06259482),
	.w8(0.06310034),
	.w9(0.073451795),
	.w10(-0.011218734),
	.w11(-0.058841117),
	.w12(0.015071797),
	.w13(-0.017841464),
	.w14(0.011094039),
	.w15(0.008163197),
	.w16(-0.04719745),
	.w17(-0.04609858),
	.w18(-0.0643243),
	.w19(0.060044125),
	.w20(-0.05405061),
	.w21(0.004496713),
	.w22(0.06512866),
	.w23(-0.0021838339),
	.w24(-0.042488005),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.027680373),
	.w1(0.02509089),
	.w2(-0.013130013),
	.w3(-0.035974815),
	.w4(-0.017565269),
	.w5(-0.011783739),
	.w6(0.057246454),
	.w7(-0.017750584),
	.w8(0.0043538753),
	.w9(0.051564086),
	.w10(0.01664237),
	.w11(0.007093905),
	.w12(-0.011086243),
	.w13(-0.08160306),
	.w14(-0.05984144),
	.w15(0.070812166),
	.w16(0.045241),
	.w17(-0.00055242877),
	.w18(0.07478075),
	.w19(0.039340887),
	.w20(0.01319803),
	.w21(-0.009610835),
	.w22(-0.0027327877),
	.w23(-0.06428234),
	.w24(0.019094279),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.06256708),
	.w1(-0.03608418),
	.w2(0.028415352),
	.w3(0.01862259),
	.w4(-0.022650493),
	.w5(0.054233667),
	.w6(-0.02549289),
	.w7(-0.019123208),
	.w8(0.062841505),
	.w9(-0.010166243),
	.w10(0.049735494),
	.w11(0.04807707),
	.w12(-0.03878323),
	.w13(0.066284046),
	.w14(-0.022285383),
	.w15(0.044601213),
	.w16(-0.05804251),
	.w17(-0.013679035),
	.w18(0.07752017),
	.w19(-0.046109375),
	.w20(-0.037827197),
	.w21(-0.008889201),
	.w22(0.044825967),
	.w23(0.03893076),
	.w24(-0.021366443),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.032637905),
	.w1(0.031061249),
	.w2(0.07461572),
	.w3(0.041664355),
	.w4(0.02118408),
	.w5(0.07606527),
	.w6(0.016559118),
	.w7(-0.035849478),
	.w8(-0.058292776),
	.w9(-0.04976413),
	.w10(0.041489594),
	.w11(-0.07210196),
	.w12(-0.031451784),
	.w13(-0.014466068),
	.w14(-0.03382235),
	.w15(0.01458282),
	.w16(-0.012552511),
	.w17(0.0052191163),
	.w18(0.07653919),
	.w19(-0.014864816),
	.w20(0.07489512),
	.w21(0.063014895),
	.w22(0.02996776),
	.w23(-0.029059205),
	.w24(-0.020527843),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.03745002),
	.w1(-0.07843338),
	.w2(0.0021067746),
	.w3(0.048544455),
	.w4(-0.010089241),
	.w5(-0.06357358),
	.w6(-0.052369848),
	.w7(-0.06869652),
	.w8(-0.024388859),
	.w9(0.007785492),
	.w10(0.07468993),
	.w11(0.016401486),
	.w12(-0.064011715),
	.w13(0.025292663),
	.w14(-0.0759018),
	.w15(0.0058098556),
	.w16(0.058774948),
	.w17(-0.02683345),
	.w18(-0.07988971),
	.w19(0.0777144),
	.w20(0.034133267),
	.w21(-0.06484887),
	.w22(-0.05890565),
	.w23(0.010000521),
	.w24(0.037399463),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.017946789),
	.w1(-0.020953923),
	.w2(0.003396703),
	.w3(-0.047456875),
	.w4(0.046527084),
	.w5(-0.01585302),
	.w6(0.08045648),
	.w7(0.06570716),
	.w8(0.019407013),
	.w9(-0.07637194),
	.w10(-0.07757158),
	.w11(0.037876993),
	.w12(-0.012545056),
	.w13(-0.012053441),
	.w14(-0.07397847),
	.w15(0.055460308),
	.w16(0.039372995),
	.w17(-0.03803922),
	.w18(0.01670732),
	.w19(-0.028843757),
	.w20(-0.0035854725),
	.w21(-0.007852332),
	.w22(-0.06117459),
	.w23(0.011939258),
	.w24(-0.04967681),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule