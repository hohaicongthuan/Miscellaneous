module featuremap5(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.058393024),
	.w1(-0.07127947),
	.w2(0.07297034),
	.w3(-0.039839964),
	.w4(0.009093379),
	.w5(-0.082046755),
	.w6(0.021941064),
	.w7(-0.06185163),
	.w8(0.0626271),
	.w9(0.06897338),
	.w10(0.0036860881),
	.w11(-0.06048919),
	.w12(0.050356697),
	.w13(0.028401606),
	.w14(-0.06634381),
	.w15(0.014039069),
	.w16(0.06187217),
	.w17(-0.032866564),
	.w18(0.10097026),
	.w19(-0.0963859),
	.w20(0.054610018),
	.w21(-0.015189708),
	.w22(-0.085940495),
	.w23(0.012705135),
	.w24(-0.054090522),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.07298946),
	.w1(-0.01703108),
	.w2(0.023676898),
	.w3(-0.09230157),
	.w4(0.00067356776),
	.w5(0.09050067),
	.w6(0.09166917),
	.w7(0.081440926),
	.w8(-0.057747222),
	.w9(0.06597457),
	.w10(0.014583218),
	.w11(-0.050342023),
	.w12(0.013515308),
	.w13(-0.042615518),
	.w14(-0.043676645),
	.w15(0.06191707),
	.w16(0.07896075),
	.w17(-0.041479446),
	.w18(0.08239445),
	.w19(0.07581005),
	.w20(-0.021595161),
	.w21(0.055300035),
	.w22(0.05140209),
	.w23(-0.041977316),
	.w24(-0.05799761),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.056461904),
	.w1(-0.058077544),
	.w2(-0.1102135),
	.w3(-0.060196184),
	.w4(0.08889998),
	.w5(0.01830983),
	.w6(0.06912394),
	.w7(0.11020274),
	.w8(0.055222344),
	.w9(0.06954146),
	.w10(-0.07017576),
	.w11(-0.060108982),
	.w12(0.082147546),
	.w13(-0.1097425),
	.w14(-0.08761996),
	.w15(-0.022140274),
	.w16(-0.041516073),
	.w17(-0.08650845),
	.w18(0.07713073),
	.w19(0.06086254),
	.w20(0.027619349),
	.w21(-0.04943694),
	.w22(0.07145305),
	.w23(0.066404216),
	.w24(-0.07310724),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule