module featuremap11(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.007800238),
	.w1(-0.0649969),
	.w2(0.028459113),
	.w3(0.047146887),
	.w4(0.025080893),
	.w5(0.018451096),
	.w6(0.017393826),
	.w7(-0.017183254),
	.w8(0.03199009),
	.w9(0.07625273),
	.w10(-0.06729105),
	.w11(-0.024615861),
	.w12(-0.04076018),
	.w13(0.03408085),
	.w14(-0.05285229),
	.w15(-0.048867352),
	.w16(-0.075198725),
	.w17(-0.0644302),
	.w18(0.04834964),
	.w19(0.0050223265),
	.w20(0.045227043),
	.w21(0.04381352),
	.w22(0.007186966),
	.w23(-0.07846585),
	.w24(-0.01344409),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.047985505),
	.w1(-0.037050404),
	.w2(0.057475697),
	.w3(0.023279533),
	.w4(0.01382018),
	.w5(0.061327085),
	.w6(0.037713412),
	.w7(0.011819159),
	.w8(0.025671829),
	.w9(0.03486589),
	.w10(-0.026452009),
	.w11(-0.013371158),
	.w12(-0.080448404),
	.w13(-0.024173137),
	.w14(0.04409174),
	.w15(0.016920324),
	.w16(0.07863509),
	.w17(-0.057714984),
	.w18(0.07227389),
	.w19(-0.05856638),
	.w20(0.019029543),
	.w21(0.034407523),
	.w22(0.003456719),
	.w23(-0.03701595),
	.w24(-0.014743314),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.030141491),
	.w1(-0.037182536),
	.w2(-0.017100295),
	.w3(0.060230356),
	.w4(0.01860505),
	.w5(0.043187495),
	.w6(-0.033890847),
	.w7(0.016360411),
	.w8(-0.052962203),
	.w9(0.002014385),
	.w10(-0.05118939),
	.w11(-0.056700043),
	.w12(-0.019345168),
	.w13(-0.04266466),
	.w14(0.021484004),
	.w15(0.025994256),
	.w16(0.057068344),
	.w17(-0.02851941),
	.w18(0.03495343),
	.w19(-0.011025555),
	.w20(-0.019025864),
	.w21(-0.08156122),
	.w22(0.018856863),
	.w23(-0.032106206),
	.w24(-0.058321733),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.0052726013),
	.w1(0.07297953),
	.w2(-0.028822627),
	.w3(-3.9001727e-05),
	.w4(0.07664748),
	.w5(-0.038337722),
	.w6(0.07898485),
	.w7(-0.00979063),
	.w8(-0.020778585),
	.w9(0.018884836),
	.w10(-0.019788262),
	.w11(-0.025741082),
	.w12(-0.07786298),
	.w13(0.04686269),
	.w14(0.0015766255),
	.w15(0.01302205),
	.w16(0.03210062),
	.w17(-0.051000107),
	.w18(-0.03357748),
	.w19(-0.008871758),
	.w20(0.024393395),
	.w21(-0.0026064678),
	.w22(0.06594042),
	.w23(-0.02306684),
	.w24(0.00075056177),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.048861932),
	.w1(0.047645975),
	.w2(0.029677996),
	.w3(0.049780305),
	.w4(0.05611594),
	.w5(-0.014285504),
	.w6(0.06580874),
	.w7(-0.0062584872),
	.w8(0.022301093),
	.w9(0.041028637),
	.w10(-0.05148488),
	.w11(0.064029284),
	.w12(-0.013918254),
	.w13(0.020374903),
	.w14(0.035285436),
	.w15(0.07914223),
	.w16(0.057227407),
	.w17(0.046962067),
	.w18(-0.0039570155),
	.w19(-0.057067584),
	.w20(-0.071897596),
	.w21(0.013354514),
	.w22(-0.072996885),
	.w23(-0.0054063965),
	.w24(-0.038121767),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.059362583),
	.w1(-0.03896033),
	.w2(-0.015091488),
	.w3(-0.020696932),
	.w4(-0.079998985),
	.w5(-0.0036475617),
	.w6(0.08016344),
	.w7(-0.06649155),
	.w8(-0.035709687),
	.w9(0.07596011),
	.w10(0.016139511),
	.w11(-0.04084168),
	.w12(-0.0061445385),
	.w13(0.00545409),
	.w14(0.056534417),
	.w15(0.028743543),
	.w16(0.060740016),
	.w17(-0.06592686),
	.w18(0.06758335),
	.w19(0.074833564),
	.w20(0.062560685),
	.w21(0.04559549),
	.w22(-0.035243154),
	.w23(0.038969588),
	.w24(-0.010605073),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule