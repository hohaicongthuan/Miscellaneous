module featuremap6(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.017831108),
	.w1(-0.008601491),
	.w2(-0.041576415),
	.w3(-0.021546755),
	.w4(0.07773062),
	.w5(-0.012925806),
	.w6(0.016584095),
	.w7(-0.055875234),
	.w8(-0.054117274),
	.w9(-0.06136451),
	.w10(0.043066002),
	.w11(0.06515316),
	.w12(-0.056386422),
	.w13(0.08132344),
	.w14(-0.02778637),
	.w15(0.07890778),
	.w16(0.0040721423),
	.w17(-0.06410036),
	.w18(0.024525875),
	.w19(0.057916258),
	.w20(-0.025827523),
	.w21(0.036365084),
	.w22(-0.043949146),
	.w23(-0.04320046),
	.w24(0.0043623243),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.04000588),
	.w1(0.026905263),
	.w2(-0.03200171),
	.w3(-0.004307603),
	.w4(0.03893485),
	.w5(-0.03690998),
	.w6(-0.010315659),
	.w7(-0.01149598),
	.w8(-0.069645025),
	.w9(-0.0396855),
	.w10(-0.07108422),
	.w11(-0.038209416),
	.w12(0.072964765),
	.w13(-0.022783423),
	.w14(0.045898598),
	.w15(0.05830073),
	.w16(-0.021246752),
	.w17(0.059622545),
	.w18(0.0061546806),
	.w19(-0.05549641),
	.w20(0.055667173),
	.w21(-0.04098737),
	.w22(-0.020983348),
	.w23(0.0018983922),
	.w24(-0.04935196),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.077522054),
	.w1(-0.08029223),
	.w2(-0.03600921),
	.w3(-0.03529264),
	.w4(0.0016632528),
	.w5(0.06234231),
	.w6(-0.009139077),
	.w7(-0.0790486),
	.w8(0.03178231),
	.w9(-0.07900349),
	.w10(0.075962104),
	.w11(0.015247427),
	.w12(-0.06673532),
	.w13(0.022437926),
	.w14(-0.050661683),
	.w15(0.059495755),
	.w16(0.00631754),
	.w17(0.027590543),
	.w18(0.070977435),
	.w19(-0.025686506),
	.w20(-0.05327489),
	.w21(-0.050090745),
	.w22(0.01237805),
	.w23(-0.06956602),
	.w24(-0.010515126),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07259756),
	.w1(0.079863),
	.w2(0.034880497),
	.w3(-0.018362124),
	.w4(0.00994472),
	.w5(-0.02457536),
	.w6(-0.020484297),
	.w7(-0.062213447),
	.w8(0.045688026),
	.w9(-0.045382015),
	.w10(-0.050131768),
	.w11(0.05988376),
	.w12(-0.019583559),
	.w13(-0.012431885),
	.w14(-0.011747492),
	.w15(-0.056211554),
	.w16(-0.06790948),
	.w17(-0.006589355),
	.w18(-0.07613568),
	.w19(0.011251662),
	.w20(-0.059727352),
	.w21(-0.008823549),
	.w22(-0.00601524),
	.w23(0.032652836),
	.w24(-0.07770554),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.0074355765),
	.w1(-0.055786),
	.w2(0.016178932),
	.w3(0.062251594),
	.w4(0.004272923),
	.w5(-0.062098194),
	.w6(0.03036643),
	.w7(0.047262978),
	.w8(0.017667918),
	.w9(-0.0057688486),
	.w10(-0.0027735513),
	.w11(0.0695099),
	.w12(0.057980392),
	.w13(0.08051901),
	.w14(0.0802604),
	.w15(-0.006149405),
	.w16(-0.03995268),
	.w17(-0.006489266),
	.w18(-0.06358998),
	.w19(-0.06944493),
	.w20(0.07846055),
	.w21(0.017616244),
	.w22(-0.04256453),
	.w23(-0.0067001693),
	.w24(-0.00064275466),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.047268633),
	.w1(-0.03874606),
	.w2(-0.027402524),
	.w3(0.05237846),
	.w4(0.06538469),
	.w5(-0.007730547),
	.w6(-0.06863151),
	.w7(-0.05330796),
	.w8(-0.041224103),
	.w9(-0.017774383),
	.w10(0.04843962),
	.w11(-0.04346403),
	.w12(-0.06546599),
	.w13(0.019732071),
	.w14(0.010977229),
	.w15(0.03406635),
	.w16(-0.027969873),
	.w17(0.009554235),
	.w18(0.08151351),
	.w19(0.060580563),
	.w20(-0.027062876),
	.w21(0.015352324),
	.w22(-0.0036582004),
	.w23(0.0035864555),
	.w24(-0.063170545),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule