module featuremap10(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.050210103),
	.w1(0.0014713005),
	.w2(-0.045446064),
	.w3(0.023164446),
	.w4(-0.009896189),
	.w5(-0.073516764),
	.w6(0.0068559623),
	.w7(0.011241461),
	.w8(-0.0012357717),
	.w9(0.006790982),
	.w10(0.04896639),
	.w11(-0.065160565),
	.w12(-0.07941227),
	.w13(0.0027780968),
	.w14(0.07871457),
	.w15(0.0023912233),
	.w16(-0.046642248),
	.w17(-0.020743283),
	.w18(0.049771808),
	.w19(-0.02821568),
	.w20(-0.02125712),
	.w21(0.056830917),
	.w22(-0.060947288),
	.w23(0.06342545),
	.w24(-0.033240616),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07265758),
	.w1(-0.00093548663),
	.w2(-0.06648174),
	.w3(0.03276254),
	.w4(0.034608033),
	.w5(-0.024026124),
	.w6(0.06783571),
	.w7(-0.07101046),
	.w8(0.02596019),
	.w9(0.004308644),
	.w10(0.075568795),
	.w11(0.005102325),
	.w12(0.036522776),
	.w13(-0.07556498),
	.w14(-0.01267159),
	.w15(0.05767633),
	.w16(0.031111006),
	.w17(0.05560331),
	.w18(-0.044460915),
	.w19(0.02850919),
	.w20(0.005570755),
	.w21(0.06326189),
	.w22(0.008317685),
	.w23(0.040989317),
	.w24(0.019868484),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.044102933),
	.w1(-0.016385077),
	.w2(-0.0788248),
	.w3(-0.051298648),
	.w4(-0.03590128),
	.w5(0.03972345),
	.w6(-0.08038467),
	.w7(-0.0112067135),
	.w8(0.073919766),
	.w9(0.052329786),
	.w10(-0.065730006),
	.w11(0.022876473),
	.w12(-0.055496965),
	.w13(-0.025056142),
	.w14(-0.048833888),
	.w15(0.04711747),
	.w16(-0.06811311),
	.w17(0.027139176),
	.w18(-0.023412619),
	.w19(-0.06802937),
	.w20(-0.013114644),
	.w21(-0.0040032202),
	.w22(-0.048763566),
	.w23(0.042113278),
	.w24(-0.07697358),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.05518085),
	.w1(0.025157807),
	.w2(-0.06435821),
	.w3(0.07336614),
	.w4(0.08112858),
	.w5(-0.048853774),
	.w6(0.04412559),
	.w7(0.025404053),
	.w8(-0.041576054),
	.w9(0.080281794),
	.w10(0.008712443),
	.w11(0.0052983556),
	.w12(-0.0044666077),
	.w13(0.04866846),
	.w14(0.06592416),
	.w15(0.052219283),
	.w16(-0.014309643),
	.w17(0.074389696),
	.w18(0.03340035),
	.w19(0.057978448),
	.w20(-0.032229003),
	.w21(0.06003998),
	.w22(-0.020753289),
	.w23(0.014132777),
	.w24(0.049736943),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07080579),
	.w1(-0.012374108),
	.w2(0.06524633),
	.w3(-0.058783066),
	.w4(0.042813607),
	.w5(0.026239168),
	.w6(-0.020352468),
	.w7(-0.054679126),
	.w8(-0.042072974),
	.w9(-0.0034867856),
	.w10(-0.0009663999),
	.w11(-0.004631735),
	.w12(-0.03679379),
	.w13(-0.051954456),
	.w14(0.03983097),
	.w15(0.033614814),
	.w16(0.05448332),
	.w17(0.033905067),
	.w18(-0.06749058),
	.w19(0.009168316),
	.w20(-0.05381907),
	.w21(-0.0718867),
	.w22(-0.032080688),
	.w23(0.073396415),
	.w24(0.021160515),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.04401573),
	.w1(0.05928642),
	.w2(-0.07248996),
	.w3(-0.051172543),
	.w4(-0.07980958),
	.w5(-0.080845974),
	.w6(-0.011587893),
	.w7(0.015608399),
	.w8(0.040548608),
	.w9(-0.019786732),
	.w10(0.07595552),
	.w11(-0.07861442),
	.w12(-0.04634142),
	.w13(-0.07951946),
	.w14(0.057736475),
	.w15(0.0009966805),
	.w16(-0.03663685),
	.w17(-0.002896854),
	.w18(0.064567044),
	.w19(-0.025194269),
	.w20(-0.07291165),
	.w21(-0.011312934),
	.w22(-0.07481733),
	.w23(-0.04161965),
	.w24(-0.022437468),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule