module featuremap2(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.021808408),
	.w1(0.04928916),
	.w2(-0.01824032),
	.w3(-0.040658332),
	.w4(0.057173718),
	.w5(-0.019273685),
	.w6(0.0103458725),
	.w7(0.03289326),
	.w8(-0.0677516),
	.w9(-0.043222964),
	.w10(0.051369946),
	.w11(0.05197903),
	.w12(0.013444879),
	.w13(0.07346697),
	.w14(-0.0041778176),
	.w15(0.05827075),
	.w16(-0.0728997),
	.w17(0.07254563),
	.w18(0.0170461),
	.w19(-0.03297533),
	.w20(0.046817567),
	.w21(-0.061925486),
	.w22(-0.074782476),
	.w23(0.019040668),
	.w24(0.04451194),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.067518346),
	.w1(-0.019148719),
	.w2(-0.02300256),
	.w3(-0.07020005),
	.w4(-0.048387118),
	.w5(-0.00028571417),
	.w6(0.020749064),
	.w7(-0.025752585),
	.w8(-0.0033974426),
	.w9(0.081127904),
	.w10(0.020419072),
	.w11(-0.0731786),
	.w12(-0.028274344),
	.w13(-0.068591595),
	.w14(-0.038744833),
	.w15(0.050944634),
	.w16(0.04147625),
	.w17(-0.016168274),
	.w18(-0.06103233),
	.w19(0.034301158),
	.w20(-0.06293582),
	.w21(-0.017784836),
	.w22(0.0703738),
	.w23(0.007805786),
	.w24(0.030163733),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.023014843),
	.w1(0.036672544),
	.w2(0.030278761),
	.w3(-0.059286516),
	.w4(-0.03676432),
	.w5(0.07168466),
	.w6(-0.010895313),
	.w7(0.077557296),
	.w8(0.036673985),
	.w9(-0.024062594),
	.w10(-0.021325845),
	.w11(0.038042404),
	.w12(0.06504016),
	.w13(-0.06301435),
	.w14(-0.011595883),
	.w15(0.014946149),
	.w16(0.021965826),
	.w17(-0.046812642),
	.w18(0.033135243),
	.w19(0.07521577),
	.w20(0.010947406),
	.w21(0.05350191),
	.w22(-0.023910696),
	.w23(0.06988467),
	.w24(0.06284751),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.068480566),
	.w1(0.026199572),
	.w2(0.06439317),
	.w3(-0.027205236),
	.w4(0.07760052),
	.w5(-0.076090686),
	.w6(0.027635405),
	.w7(0.0046987007),
	.w8(0.028131964),
	.w9(-0.034707904),
	.w10(-0.028935192),
	.w11(-0.058002632),
	.w12(0.015547069),
	.w13(-0.014262718),
	.w14(-0.0027499478),
	.w15(0.06924968),
	.w16(0.051191628),
	.w17(-0.043253236),
	.w18(0.0654174),
	.w19(0.014947414),
	.w20(-0.021876201),
	.w21(0.04314605),
	.w22(0.006980754),
	.w23(-0.08146823),
	.w24(-0.0016301203),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.037491065),
	.w1(-0.02681663),
	.w2(-0.05763368),
	.w3(-0.034438077),
	.w4(-0.071868025),
	.w5(0.0047036256),
	.w6(-0.03565997),
	.w7(0.048606936),
	.w8(-0.0555643),
	.w9(-0.04617125),
	.w10(0.06601194),
	.w11(-0.032657634),
	.w12(0.047945287),
	.w13(0.04774993),
	.w14(0.06680926),
	.w15(0.0498634),
	.w16(-0.04730811),
	.w17(0.038900673),
	.w18(-0.037403893),
	.w19(-0.0568885),
	.w20(0.05859134),
	.w21(0.044012498),
	.w22(0.048824206),
	.w23(0.036741797),
	.w24(-0.05962811),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.037871853),
	.w1(-0.031600207),
	.w2(0.0018182572),
	.w3(0.009722896),
	.w4(0.011832211),
	.w5(0.05487026),
	.w6(0.023638735),
	.w7(-0.06849587),
	.w8(-0.0050093224),
	.w9(-0.047159977),
	.w10(0.047545314),
	.w11(0.0034566508),
	.w12(0.004219331),
	.w13(-0.0047535775),
	.w14(0.0732448),
	.w15(-0.062825166),
	.w16(0.058250863),
	.w17(-0.07057459),
	.w18(-0.008617464),
	.w19(-0.061809286),
	.w20(-0.021379953),
	.w21(-0.0515851),
	.w22(-0.009026403),
	.w23(0.07220546),
	.w24(0.053966973),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule