module featuremap0(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.07135645),
	.w1(-0.04893036),
	.w2(-0.0495103),
	.w3(0.02537423),
	.w4(0.0063254824),
	.w5(-0.031082993),
	.w6(0.077751875),
	.w7(0.010892928),
	.w8(0.008886437),
	.w9(-0.030188758),
	.w10(-0.075471394),
	.w11(0.022980426),
	.w12(0.08101609),
	.w13(0.08078232),
	.w14(0.042373627),
	.w15(0.01180998),
	.w16(-0.0026716914),
	.w17(-0.058708984),
	.w18(0.02854611),
	.w19(-0.0393251),
	.w20(-0.010156294),
	.w21(0.05615498),
	.w22(0.038001474),
	.w23(-0.040470157),
	.w24(0.026625585),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07048175),
	.w1(0.00039267447),
	.w2(-0.010628423),
	.w3(-0.025440533),
	.w4(0.07130053),
	.w5(-0.043205637),
	.w6(-0.06965281),
	.w7(0.03704616),
	.w8(-0.06232331),
	.w9(0.03972953),
	.w10(-0.0552087),
	.w11(0.009361524),
	.w12(0.03059136),
	.w13(0.06253855),
	.w14(0.061562177),
	.w15(0.07837431),
	.w16(-0.06094719),
	.w17(-0.016154306),
	.w18(0.007630556),
	.w19(0.012625415),
	.w20(0.007633028),
	.w21(-0.06668971),
	.w22(-0.026793174),
	.w23(-0.08072282),
	.w24(0.007417307),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.04484555),
	.w1(0.07399073),
	.w2(-0.013502024),
	.w3(-0.0023288713),
	.w4(0.016259875),
	.w5(-0.010757653),
	.w6(0.06483176),
	.w7(0.009904005),
	.w8(-0.058807265),
	.w9(0.0048643434),
	.w10(0.06162082),
	.w11(-0.008931415),
	.w12(-0.013780935),
	.w13(-0.0075789103),
	.w14(-0.0126834065),
	.w15(-0.041457463),
	.w16(0.0338787),
	.w17(-0.02109135),
	.w18(-0.030832758),
	.w19(0.07698133),
	.w20(0.039449688),
	.w21(0.0035380903),
	.w22(0.050136957),
	.w23(-0.063555345),
	.w24(0.04175627),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.05290249),
	.w1(-0.036819313),
	.w2(0.059819244),
	.w3(-0.08144434),
	.w4(-0.08110631),
	.w5(-0.027468925),
	.w6(0.064483896),
	.w7(-0.07965221),
	.w8(-0.009950599),
	.w9(-0.009394286),
	.w10(-0.05336969),
	.w11(-0.04185548),
	.w12(0.0015688777),
	.w13(-0.02306833),
	.w14(0.06417856),
	.w15(0.062095694),
	.w16(0.04366864),
	.w17(-0.07027701),
	.w18(0.0095337955),
	.w19(0.014054541),
	.w20(0.0370386),
	.w21(-0.008989611),
	.w22(0.050932147),
	.w23(0.041390557),
	.w24(-0.060732823),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.063024685),
	.w1(-0.04283358),
	.w2(0.06505738),
	.w3(-0.02818941),
	.w4(-0.018932724),
	.w5(0.04984408),
	.w6(0.06375798),
	.w7(0.012248206),
	.w8(0.01224732),
	.w9(-0.020026146),
	.w10(-0.045187175),
	.w11(-0.024303019),
	.w12(-0.019214272),
	.w13(0.023146644),
	.w14(0.08116728),
	.w15(0.04462839),
	.w16(-0.05535846),
	.w17(0.04644409),
	.w18(0.040030118),
	.w19(-0.06188432),
	.w20(0.02267073),
	.w21(0.050150614),
	.w22(0.046947137),
	.w23(0.04619473),
	.w24(0.05562092),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.0701523),
	.w1(-0.08018797),
	.w2(-0.07932805),
	.w3(0.016130071),
	.w4(0.047517624),
	.w5(-0.017392142),
	.w6(0.015956767),
	.w7(-0.0599739),
	.w8(-0.009324459),
	.w9(0.050328977),
	.w10(0.026752926),
	.w11(-0.0040377444),
	.w12(-0.059956603),
	.w13(0.03208348),
	.w14(0.020622948),
	.w15(0.010300495),
	.w16(-0.072985284),
	.w17(-0.04735599),
	.w18(0.07168059),
	.w19(0.07305857),
	.w20(0.06325136),
	.w21(-0.0574606),
	.w22(-0.041202478),
	.w23(0.05272976),
	.w24(-0.032549124),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule