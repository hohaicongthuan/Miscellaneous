module featuremap4(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(-0.009623926),
	.w1(-0.0059584165),
	.w2(0.006201333),
	.w3(-0.061589077),
	.w4(0.052861694),
	.w5(0.056883972),
	.w6(0.045203343),
	.w7(-0.044682108),
	.w8(-0.016932083),
	.w9(-0.034847803),
	.w10(0.07684402),
	.w11(-0.01371392),
	.w12(-0.02185876),
	.w13(-0.0789458),
	.w14(-0.06577628),
	.w15(0.0144090885),
	.w16(-0.0218879),
	.w17(-0.059427682),
	.w18(-0.06432867),
	.w19(-0.0012716783),
	.w20(-0.044590976),
	.w21(0.07179423),
	.w22(-0.0759857),
	.w23(-0.045313787),
	.w24(0.04798173),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.07941868),
	.w1(0.040707182),
	.w2(-0.056096707),
	.w3(0.059979994),
	.w4(0.020255037),
	.w5(-0.049671166),
	.w6(-0.05124493),
	.w7(-0.068510555),
	.w8(0.03305719),
	.w9(0.05096522),
	.w10(-0.064675964),
	.w11(-0.0241142),
	.w12(0.07042502),
	.w13(-0.012262281),
	.w14(0.017767442),
	.w15(-0.08026842),
	.w16(-0.0224031),
	.w17(0.07569898),
	.w18(0.023826707),
	.w19(-0.068229444),
	.w20(-0.046890695),
	.w21(0.04464337),
	.w22(-0.06646009),
	.w23(0.054811947),
	.w24(0.070169255),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.0021043315),
	.w1(0.07633502),
	.w2(0.02663631),
	.w3(0.07506819),
	.w4(-0.06979765),
	.w5(-0.02693829),
	.w6(-0.04147838),
	.w7(-0.045025017),
	.w8(0.025022328),
	.w9(-0.028235722),
	.w10(0.019595822),
	.w11(0.01940423),
	.w12(-0.030753898),
	.w13(-0.028322505),
	.w14(-0.077477515),
	.w15(0.015563879),
	.w16(-0.010147125),
	.w17(-0.07105083),
	.w18(-0.07815101),
	.w19(-0.03341963),
	.w20(-0.07306627),
	.w21(0.04422024),
	.w22(-0.050240763),
	.w23(-0.05673908),
	.w24(-0.07979624),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.06206729),
	.w1(0.075921774),
	.w2(-0.0034259032),
	.w3(-0.05716709),
	.w4(-0.07706931),
	.w5(-0.0048034904),
	.w6(0.02499196),
	.w7(0.043436047),
	.w8(0.014956291),
	.w9(-0.066853374),
	.w10(-0.07833323),
	.w11(0.0014539555),
	.w12(0.075577654),
	.w13(0.042563256),
	.w14(0.07716051),
	.w15(0.04297557),
	.w16(0.064381406),
	.w17(-0.07236373),
	.w18(-0.07442691),
	.w19(-0.04986857),
	.w20(0.071600884),
	.w21(0.032079276),
	.w22(0.00028177214),
	.w23(-0.058579978),
	.w24(-3.145834e-05),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.04901902),
	.w1(-0.013763492),
	.w2(0.07843761),
	.w3(0.07041773),
	.w4(-0.022750797),
	.w5(0.06949284),
	.w6(-0.07013603),
	.w7(0.000839856),
	.w8(0.024649598),
	.w9(0.04446485),
	.w10(-0.002141844),
	.w11(0.0697848),
	.w12(0.06075373),
	.w13(-0.06911578),
	.w14(0.053690854),
	.w15(0.07061321),
	.w16(0.02972466),
	.w17(-0.053200193),
	.w18(-0.04872316),
	.w19(-0.04549437),
	.w20(-0.0036922088),
	.w21(0.06631375),
	.w22(0.046504024),
	.w23(0.055228915),
	.w24(0.047186464),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.023641393),
	.w1(-0.03630492),
	.w2(-0.05305166),
	.w3(-0.035635266),
	.w4(0.056688264),
	.w5(0.076927036),
	.w6(0.05798454),
	.w7(-0.036933154),
	.w8(-0.04079972),
	.w9(0.021811046),
	.w10(0.032509822),
	.w11(0.07563058),
	.w12(-0.045427103),
	.w13(0.032534905),
	.w14(0.023490222),
	.w15(-0.0316176),
	.w16(-0.039922953),
	.w17(0.03964093),
	.w18(-0.068429105),
	.w19(-0.029498134),
	.w20(-0.06592156),
	.w21(-0.020738173),
	.w22(0.030287318),
	.w23(0.05121124),
	.w24(-0.0043499335),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule