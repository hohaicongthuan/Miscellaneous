module featuremap7(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.0006421804),
	.w1(0.08081481),
	.w2(-0.016735507),
	.w3(-0.04730779),
	.w4(0.030053608),
	.w5(-0.019409573),
	.w6(0.037097562),
	.w7(0.048241828),
	.w8(-0.067002825),
	.w9(0.04081675),
	.w10(0.01147299),
	.w11(0.039694734),
	.w12(0.0063514123),
	.w13(-0.05288385),
	.w14(-0.06708327),
	.w15(-0.0604211),
	.w16(0.03916987),
	.w17(-0.013378877),
	.w18(0.023385901),
	.w19(-0.032614738),
	.w20(0.045507364),
	.w21(-0.06933907),
	.w22(0.06482454),
	.w23(0.012991117),
	.w24(-0.051066283),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.0081437295),
	.w1(-0.075045764),
	.w2(-0.038334113),
	.w3(0.07327489),
	.w4(0.045772716),
	.w5(-0.008398988),
	.w6(0.030725028),
	.w7(-0.042839225),
	.w8(0.0184437),
	.w9(-0.07140306),
	.w10(-0.07715281),
	.w11(-0.058019094),
	.w12(-0.061298996),
	.w13(-0.05722182),
	.w14(-0.07069173),
	.w15(-0.07153647),
	.w16(-0.06656711),
	.w17(-0.024448972),
	.w18(-0.064036),
	.w19(-0.06126844),
	.w20(0.061270796),
	.w21(0.02701309),
	.w22(0.04302527),
	.w23(0.01992993),
	.w24(0.077959515),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.06265529),
	.w1(-0.059735615),
	.w2(-0.020379672),
	.w3(-0.050056696),
	.w4(0.072240755),
	.w5(-0.08028061),
	.w6(-0.027557168),
	.w7(0.032162573),
	.w8(-0.06831852),
	.w9(0.0022830658),
	.w10(0.07496275),
	.w11(0.063700914),
	.w12(0.019201085),
	.w13(0.06389879),
	.w14(-0.074054755),
	.w15(-0.045634452),
	.w16(0.055616695),
	.w17(-0.02139251),
	.w18(0.011372318),
	.w19(0.016761145),
	.w20(0.036317237),
	.w21(0.056843095),
	.w22(-0.048736855),
	.w23(-0.010161697),
	.w24(-0.048012946),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.049211554),
	.w1(0.027461313),
	.w2(0.037361484),
	.w3(-0.027210414),
	.w4(0.035182294),
	.w5(-0.03734338),
	.w6(-0.005618137),
	.w7(-0.053948984),
	.w8(0.02034213),
	.w9(0.0052361107),
	.w10(0.025592588),
	.w11(0.030549778),
	.w12(0.04275877),
	.w13(0.034876682),
	.w14(-0.04620782),
	.w15(-0.06090957),
	.w16(0.02801124),
	.w17(0.059533462),
	.w18(0.025456592),
	.w19(-0.014718514),
	.w20(-0.0543259),
	.w21(0.020252846),
	.w22(0.017994804),
	.w23(0.080778174),
	.w24(0.004451774),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.043309554),
	.w1(-0.07339305),
	.w2(-0.00036182933),
	.w3(0.050209843),
	.w4(0.009452531),
	.w5(0.07073233),
	.w6(0.06366746),
	.w7(-0.07719621),
	.w8(-0.017322792),
	.w9(-0.010044195),
	.w10(-0.04467621),
	.w11(0.07138269),
	.w12(0.06114757),
	.w13(0.051855896),
	.w14(0.009168335),
	.w15(0.021797847),
	.w16(-0.033987977),
	.w17(-0.056478754),
	.w18(0.045456927),
	.w19(0.07446401),
	.w20(-0.010090701),
	.w21(-0.024270734),
	.w22(-0.075571254),
	.w23(-0.015206439),
	.w24(-0.014370798),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.042963725),
	.w1(0.006314513),
	.w2(0.0051575718),
	.w3(-0.06731306),
	.w4(-0.042343408),
	.w5(-0.04589782),
	.w6(-0.08146248),
	.w7(-0.021152368),
	.w8(-0.060558848),
	.w9(0.03832327),
	.w10(0.07469641),
	.w11(-0.059331533),
	.w12(-0.06953635),
	.w13(0.056806993),
	.w14(-0.04259373),
	.w15(-0.03326084),
	.w16(0.012165706),
	.w17(-0.06347715),
	.w18(-0.045926504),
	.w19(0.06833245),
	.w20(0.013294147),
	.w21(-0.027679244),
	.w22(0.038201854),
	.w23(0.035352472),
	.w24(-0.02106504),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule