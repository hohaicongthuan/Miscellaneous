module featuremap8(
	input clk,
	input rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_WIDTH = 24;
conv2d5x5 #(
	.w0(0.0022802334),
	.w1(-0.049570777),
	.w2(0.06739196),
	.w3(0.05617329),
	.w4(-0.039704595),
	.w5(0.018824255),
	.w6(0.002989039),
	.w7(0.023105461),
	.w8(0.04379744),
	.w9(-0.020346053),
	.w10(-0.07852012),
	.w11(0.0115242265),
	.w12(0.0055049667),
	.w13(0.06658185),
	.w14(0.0067289514),
	.w15(-0.05418718),
	.w16(-0.022648644),
	.w17(0.0010303872),
	.w18(-0.024287952),
	.w19(0.0465374),
	.w20(0.040554825),
	.w21(0.041441157),
	.w22(-0.08081236),
	.w23(-0.048634548),
	.w24(-0.047434032),
)
conv2d5x5_inst0(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.027247606),
	.w1(-0.001145144),
	.w2(0.075332455),
	.w3(-0.0779632),
	.w4(0.045017473),
	.w5(-0.0015697927),
	.w6(0.07485243),
	.w7(0.011493002),
	.w8(-0.05012518),
	.w9(0.02402845),
	.w10(-0.04013078),
	.w11(-0.027577968),
	.w12(-0.06423753),
	.w13(0.03539052),
	.w14(-0.0005890166),
	.w15(-0.022604775),
	.w16(-0.014318053),
	.w17(-0.064628296),
	.w18(-0.02778456),
	.w19(-0.006219651),
	.w20(-0.061591074),
	.w21(0.045858875),
	.w22(-0.015013027),
	.w23(0.043071903),
	.w24(0.03330139),
)
conv2d5x5_inst1(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.029289274),
	.w1(0.02410914),
	.w2(-0.079203345),
	.w3(-0.028679408),
	.w4(0.010631236),
	.w5(0.002083278),
	.w6(0.012709628),
	.w7(-0.077109344),
	.w8(0.0782071),
	.w9(-0.06889989),
	.w10(-0.009592234),
	.w11(-0.04735344),
	.w12(0.008347703),
	.w13(0.047930513),
	.w14(-0.059400827),
	.w15(0.058182634),
	.w16(-0.038624372),
	.w17(0.038428847),
	.w18(-0.042938225),
	.w19(0.07759006),
	.w20(0.009479727),
	.w21(0.07403809),
	.w22(0.03476542),
	.w23(0.061715495),
	.w24(-0.037604973),
)
conv2d5x5_inst2(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.07651318),
	.w1(0.03619508),
	.w2(0.021316482),
	.w3(-0.079673395),
	.w4(0.07435407),
	.w5(-0.010781763),
	.w6(0.015696302),
	.w7(0.048159286),
	.w8(-0.064090006),
	.w9(-0.0019197083),
	.w10(0.035658665),
	.w11(-0.052051857),
	.w12(-0.019870061),
	.w13(-0.000698858),
	.w14(0.047056686),
	.w15(-0.010348569),
	.w16(-0.047244318),
	.w17(-0.057999898),
	.w18(-0.021844335),
	.w19(-0.075242065),
	.w20(-0.047811046),
	.w21(-0.023564285),
	.w22(-0.076743335),
	.w23(-0.045540914),
	.w24(0.077407956),
)
conv2d5x5_inst3(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(0.0291401),
	.w1(-0.043568872),
	.w2(-0.029068423),
	.w3(-0.067567915),
	.w4(0.042209804),
	.w5(-0.027327634),
	.w6(0.048819035),
	.w7(-0.0032434894),
	.w8(0.06787324),
	.w9(0.015121574),
	.w10(-0.025079278),
	.w11(-0.03317665),
	.w12(0.036079224),
	.w13(-0.027978994),
	.w14(-0.029956557),
	.w15(-0.020108782),
	.w16(-0.041526735),
	.w17(0.06178943),
	.w18(-0.043207984),
	.w19(-0.027084349),
	.w20(-0.040033877),
	.w21(-0.070671916),
	.w22(0.024963751),
	.w23(0.053973008),
	.w24(-0.064934105),
)
conv2d5x5_inst4(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

conv2d5x5 #(
	.w0(-0.048360847),
	.w1(-0.06584902),
	.w2(0.061016046),
	.w3(-0.061970357),
	.w4(-0.04200522),
	.w5(-0.061227705),
	.w6(0.02501566),
	.w7(-0.006304351),
	.w8(0.03503091),
	.w9(0.042126488),
	.w10(-0.05420847),
	.w11(0.042145777),
	.w12(0.06539105),
	.w13(-0.06910311),
	.w14(-0.017162755),
	.w15(-0.004479037),
	.w16(-0.05851764),
	.w17(-0.0056815404),
	.w18(-0.028579388),
	.w19(-0.039357647),
	.w20(-0.008658092),
	.w21(0.029959993),
	.w22(-0.04941134),
	.w23(-0.016221438),
	.w24(0.06644922),
)
conv2d5x5_inst5(
	.clk(clk),
	.rst(rst),
	.data_in(data_in),
	.valid_in(valid_in),
	.data_out(data_out),
	.valid_out(valid_out)
);

endmodule